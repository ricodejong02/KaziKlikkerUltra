q1jvfhvv.lea
